`timescale 1ns / 1ps
`default_nettype none

module sin_lut #(
    parameter integer SIN_WIDTH = 16,         // Width of sine values
    parameter integer ANGLE_WIDTH = 7        // Width of input angle (e.g., 0-127 for 128 entries)
)(
    input  logic [ANGLE_WIDTH-1:0] angle,     // Input angle (e.g., 0-127 for 0° to 180°)
    output logic [SIN_WIDTH-1:0] sin_value // Output sine value
);

    // LUT size: 2^ANGLE_WIDTH
    localparam integer SIN_LUT_SIZE = 1 << ANGLE_WIDTH;

    // Sine LUT array
    logic [SIN_WIDTH-1:0] sine_table [0:SIN_LUT_SIZE-1];

    // Precomputed sine values (16-bit fixed-point, scaled to [-32768, 32767])
    initial begin
        sine_table[0] = 0;       // sin(0.0°)
        sine_table[1] = 1608;       // sin(1.4°)
        sine_table[2] = 3215;       // sin(2.8°)
        sine_table[3] = 4821;       // sin(4.2°)
        sine_table[4] = 6423;       // sin(5.6°)
        sine_table[5] = 8022;       // sin(7.0°)
        sine_table[6] = 9615;       // sin(8.4°)
        sine_table[7] = 11203;       // sin(9.8°)
        sine_table[8] = 12785;       // sin(11.2°)
        sine_table[9] = 14358;       // sin(12.7°)
        sine_table[10] = 15923;       // sin(14.1°)
        sine_table[11] = 17479;       // sin(15.5°)
        sine_table[12] = 19023;       // sin(16.9°)
        sine_table[13] = 20557;       // sin(18.3°)
        sine_table[14] = 22078;       // sin(19.7°)
        sine_table[15] = 23585;       // sin(21.1°)
        sine_table[16] = 25079;       // sin(22.5°)
        sine_table[17] = 26557;       // sin(23.9°)
        sine_table[18] = 28019;       // sin(25.3°)
        sine_table[19] = 29465;       // sin(26.7°)
        sine_table[20] = 30892;       // sin(28.1°)
        sine_table[21] = 32302;       // sin(29.5°)
        sine_table[22] = 33691;       // sin(30.9°)
        sine_table[23] = 35061;       // sin(32.3°)
        sine_table[24] = 36409;       // sin(33.8°)
        sine_table[25] = 37735;       // sin(35.2°)
        sine_table[26] = 39039;       // sin(36.6°)
        sine_table[27] = 40319;       // sin(38.0°)
        sine_table[28] = 41574;       // sin(39.4°)
        sine_table[29] = 42805;       // sin(40.8°)
        sine_table[30] = 44010;       // sin(42.2°)
        sine_table[31] = 45189;       // sin(43.6°)
        sine_table[32] = 46340;       // sin(45.0°)
        sine_table[33] = 47463;       // sin(46.4°)
        sine_table[34] = 48558;       // sin(47.8°)
        sine_table[35] = 49623;       // sin(49.2°)
        sine_table[36] = 50659;       // sin(50.6°)
        sine_table[37] = 51664;       // sin(52.0°)
        sine_table[38] = 52638;       // sin(53.4°)
        sine_table[39] = 53580;       // sin(54.8°)
        sine_table[40] = 54490;       // sin(56.2°)
        sine_table[41] = 55367;       // sin(57.7°)
        sine_table[42] = 56211;       // sin(59.1°)
        sine_table[43] = 57021;       // sin(60.5°)
        sine_table[44] = 57796;       // sin(61.9°)
        sine_table[45] = 58537;       // sin(63.3°)
        sine_table[46] = 59242;       // sin(64.7°)
        sine_table[47] = 59912;       // sin(66.1°)
        sine_table[48] = 60546;       // sin(67.5°)
        sine_table[49] = 61143;       // sin(68.9°)
        sine_table[50] = 61704;       // sin(70.3°)
        sine_table[51] = 62227;       // sin(71.7°)
        sine_table[52] = 62713;       // sin(73.1°)
        sine_table[53] = 63161;       // sin(74.5°)
        sine_table[54] = 63570;       // sin(75.9°)
        sine_table[55] = 63942;       // sin(77.3°)
        sine_table[56] = 64275;       // sin(78.8°)
        sine_table[57] = 64570;       // sin(80.2°)
        sine_table[58] = 64825;       // sin(81.6°)
        sine_table[59] = 65042;       // sin(83.0°)
        sine_table[60] = 65219;       // sin(84.4°)
        sine_table[61] = 65357;       // sin(85.8°)
        sine_table[62] = 65456;       // sin(87.2°)
        sine_table[63] = 65515;       // sin(88.6°)
        sine_table[64] = 65535;       // sin(90.0°)
        sine_table[65] = 65515;       // sin(91.4°)
        sine_table[66] = 65456;       // sin(92.8°)
        sine_table[67] = 65357;       // sin(94.2°)
        sine_table[68] = 65219;       // sin(95.6°)
        sine_table[69] = 65042;       // sin(97.0°)
        sine_table[70] = 64825;       // sin(98.4°)
        sine_table[71] = 64570;       // sin(99.8°)
        sine_table[72] = 64275;       // sin(101.2°)
        sine_table[73] = 63942;       // sin(102.7°)
        sine_table[74] = 63570;       // sin(104.1°)
        sine_table[75] = 63161;       // sin(105.5°)
        sine_table[76] = 62713;       // sin(106.9°)
        sine_table[77] = 62227;       // sin(108.3°)
        sine_table[78] = 61704;       // sin(109.7°)
        sine_table[79] = 61143;       // sin(111.1°)
        sine_table[80] = 60546;       // sin(112.5°)
        sine_table[81] = 59912;       // sin(113.9°)
        sine_table[82] = 59242;       // sin(115.3°)
        sine_table[83] = 58537;       // sin(116.7°)
        sine_table[84] = 57796;       // sin(118.1°)
        sine_table[85] = 57021;       // sin(119.5°)
        sine_table[86] = 56211;       // sin(120.9°)
        sine_table[87] = 55367;       // sin(122.3°)
        sine_table[88] = 54490;       // sin(123.8°)
        sine_table[89] = 53580;       // sin(125.2°)
        sine_table[90] = 52638;       // sin(126.6°)
        sine_table[91] = 51664;       // sin(128.0°)
        sine_table[92] = 50659;       // sin(129.4°)
        sine_table[93] = 49623;       // sin(130.8°)
        sine_table[94] = 48558;       // sin(132.2°)
        sine_table[95] = 47463;       // sin(133.6°)
        sine_table[96] = 46340;       // sin(135.0°)
        sine_table[97] = 45189;       // sin(136.4°)
        sine_table[98] = 44010;       // sin(137.8°)
        sine_table[99] = 42805;       // sin(139.2°)
        sine_table[100] = 41574;       // sin(140.6°)
        sine_table[101] = 40319;       // sin(142.0°)
        sine_table[102] = 39039;       // sin(143.4°)
        sine_table[103] = 37735;       // sin(144.8°)
        sine_table[104] = 36409;       // sin(146.2°)
        sine_table[105] = 35061;       // sin(147.7°)
        sine_table[106] = 33691;       // sin(149.1°)
        sine_table[107] = 32302;       // sin(150.5°)
        sine_table[108] = 30892;       // sin(151.9°)
        sine_table[109] = 29465;       // sin(153.3°)
        sine_table[110] = 28019;       // sin(154.7°)
        sine_table[111] = 26557;       // sin(156.1°)
        sine_table[112] = 25079;       // sin(157.5°)
        sine_table[113] = 23585;       // sin(158.9°)
        sine_table[114] = 22078;       // sin(160.3°)
        sine_table[115] = 20557;       // sin(161.7°)
        sine_table[116] = 19023;       // sin(163.1°)
        sine_table[117] = 17479;       // sin(164.5°)
        sine_table[118] = 15923;       // sin(165.9°)
        sine_table[119] = 14358;       // sin(167.3°)
        sine_table[120] = 12785;       // sin(168.8°)
        sine_table[121] = 11203;       // sin(170.2°)
        sine_table[122] = 9615;       // sin(171.6°)
        sine_table[123] = 8022;       // sin(173.0°)
        sine_table[124] = 6423;       // sin(174.4°)
        sine_table[125] = 4821;       // sin(175.8°)
        sine_table[126] = 3215;       // sin(177.2°)
        sine_table[127] = 1608;       // sin(178.6°)
    end

    // Map input angle to LUT value
    assign sin_value = sine_table[angle];

endmodule

`default_nettype wire