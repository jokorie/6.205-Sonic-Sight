`timescale 1ns / 1ps
`default_nettype none

module sin_lut #(
    parameter integer SIN_WIDTH = 16,         // Width of sine values
    parameter integer ANGLE_WIDTH = 7        // Width of input angle (e.g., 0-127 for 128 entries)
)(
    input  logic signed [ANGLE_WIDTH-1:0] angle,     // Input angle (e.g., 0-127 for 0° to 180°)
    output logic [SIN_WIDTH-1:0] sin_value, // Output sine value
    output logic sign_bit  // high is negative output
);

    // LUT size: 2^ANGLE_WIDTH
    localparam integer SIN_LUT_SIZE = 1 << ANGLE_WIDTH;

    // Sine LUT array
    logic [SIN_WIDTH-1:0] cos_table [0:SIN_LUT_SIZE-1];

    // Precomputed sine values (16-bit fixed-point, scaled to [-32768, 32767])
    initial begin
        cos_table[0] = 32767;       // cos(0.0°)
        cos_table[1] = 32757;       // cos(1.4°)
        cos_table[2] = 32727;       // cos(2.8°)
        cos_table[3] = 32678;       // cos(4.2°)
        cos_table[4] = 32609;       // cos(5.6°)
        cos_table[5] = 32520;       // cos(7.0°)
        cos_table[6] = 32412;       // cos(8.4°)
        cos_table[7] = 32284;       // cos(9.8°)
        cos_table[8] = 32137;       // cos(11.2°)
        cos_table[9] = 31970;       // cos(12.7°)
        cos_table[10] = 31785;       // cos(14.1°)
        cos_table[11] = 31580;       // cos(15.5°)
        cos_table[12] = 31356;       // cos(16.9°)
        cos_table[13] = 31113;       // cos(18.3°)
        cos_table[14] = 30851;       // cos(19.7°)
        cos_table[15] = 30571;       // cos(21.1°)
        cos_table[16] = 30272;       // cos(22.5°)
        cos_table[17] = 29955;       // cos(23.9°)
        cos_table[18] = 29621;       // cos(25.3°)
        cos_table[19] = 29268;       // cos(26.7°)
        cos_table[20] = 28897;       // cos(28.1°)
        cos_table[21] = 28510;       // cos(29.5°)
        cos_table[22] = 28105;       // cos(30.9°)
        cos_table[23] = 27683;       // cos(32.3°)
        cos_table[24] = 27244;       // cos(33.8°)
        cos_table[25] = 26789;       // cos(35.2°)
        cos_table[26] = 26318;       // cos(36.6°)
        cos_table[27] = 25831;       // cos(38.0°)
        cos_table[28] = 25329;       // cos(39.4°)
        cos_table[29] = 24811;       // cos(40.8°)
        cos_table[30] = 24278;       // cos(42.2°)
        cos_table[31] = 23731;       // cos(43.6°)
        cos_table[32] = 23169;       // cos(45.0°)
        cos_table[33] = 22594;       // cos(46.4°)
        cos_table[34] = 22004;       // cos(47.8°)
        cos_table[35] = 21402;       // cos(49.2°)
        cos_table[36] = 20787;       // cos(50.6°)
        cos_table[37] = 20159;       // cos(52.0°)
        cos_table[38] = 19519;       // cos(53.4°)
        cos_table[39] = 18867;       // cos(54.8°)
        cos_table[40] = 18204;       // cos(56.2°)
        cos_table[41] = 17530;       // cos(57.7°)
        cos_table[42] = 16845;       // cos(59.1°)
        cos_table[43] = 16150;       // cos(60.5°)
        cos_table[44] = 15446;       // cos(61.9°)
        cos_table[45] = 14732;       // cos(63.3°)
        cos_table[46] = 14009;       // cos(64.7°)
        cos_table[47] = 13278;       // cos(66.1°)
        cos_table[48] = 12539;       // cos(67.5°)
        cos_table[49] = 11792;       // cos(68.9°)
        cos_table[50] = 11038;       // cos(70.3°)
        cos_table[51] = 10278;       // cos(71.7°)
        cos_table[52] = 9511;       // cos(73.1°)
        cos_table[53] = 8739;       // cos(74.5°)
        cos_table[54] = 7961;       // cos(75.9°)
        cos_table[55] = 7179;       // cos(77.3°)
        cos_table[56] = 6392;       // cos(78.8°)
        cos_table[57] = 5601;       // cos(80.2°)
        cos_table[58] = 4807;       // cos(81.6°)
        cos_table[59] = 4011;       // cos(83.0°)
        cos_table[60] = 3211;       // cos(84.4°)
        cos_table[61] = 2410;       // cos(85.8°)
        cos_table[62] = 1607;       // cos(87.2°)
        cos_table[63] = 804;       // cos(88.6°)
        cos_table[64] = 0;       // cos(90.0°)

        // TURNING POINT. BEYOND VALUES ARE ACTUALLY NEGATIVE
        cos_table[65] = 804;       // cos(91.4°)
        cos_table[66] = 1607;       // cos(92.8°)
        cos_table[67] = 2410;       // cos(94.2°)
        cos_table[68] = 3211;       // cos(95.6°)
        cos_table[69] = 4011;       // cos(97.0°)
        cos_table[70] = 4807;       // cos(98.4°)
        cos_table[71] = 5601;       // cos(99.8°)
        cos_table[72] = 6392;       // cos(101.2°)
        cos_table[73] = 7179;       // cos(102.7°)
        cos_table[74] = 7961;       // cos(104.1°)
        cos_table[75] = 8739;       // cos(105.5°)
        cos_table[76] = 9511;       // cos(106.9°)
        cos_table[77] = 10278;       // cos(108.3°)
        cos_table[78] = 11038;       // cos(109.7°)
        cos_table[79] = 11792;       // cos(111.1°)
        cos_table[80] = 12539;       // cos(112.5°)
        cos_table[81] = 13278;       // cos(113.9°)
        cos_table[82] = 14009;       // cos(115.3°)
        cos_table[83] = 14732;       // cos(116.7°)
        cos_table[84] = 15446;       // cos(118.1°)
        cos_table[85] = 16150;       // cos(119.5°)
        cos_table[86] = 16845;       // cos(120.9°)
        cos_table[87] = 17530;       // cos(122.3°)
        cos_table[88] = 18204;       // cos(123.8°)
        cos_table[89] = 18867;       // cos(125.2°)
        cos_table[90] = 19519;       // cos(126.6°)
        cos_table[91] = 20159;       // cos(128.0°)
        cos_table[92] = 20787;       // cos(129.4°)
        cos_table[93] = 21402;       // cos(130.8°)
        cos_table[94] = 22004;       // cos(132.2°)
        cos_table[95] = 22594;       // cos(133.6°)
        cos_table[96] = 23169;       // cos(135.0°)
        cos_table[97] = 23731;       // cos(136.4°)
        cos_table[98] = 24278;       // cos(137.8°)
        cos_table[99] = 24811;       // cos(139.2°)
        cos_table[100] = 25329;       // cos(140.6°)
        cos_table[101] = 25831;       // cos(142.0°)
        cos_table[102] = 26318;       // cos(143.4°)
        cos_table[103] = 26789;       // cos(144.8°)
        cos_table[104] = 27244;       // cos(146.2°)
        cos_table[105] = 27683;       // cos(147.7°)
        cos_table[106] = 28105;       // cos(149.1°)
        cos_table[107] = 28510;       // cos(150.5°)
        cos_table[108] = 28897;       // cos(151.9°)
        cos_table[109] = 29268;       // cos(153.3°)
        cos_table[110] = 29621;       // cos(154.7°)
        cos_table[111] = 29955;       // cos(156.1°)
        cos_table[112] = 30272;       // cos(157.5°)
        cos_table[113] = 30571;       // cos(158.9°)
        cos_table[114] = 30851;       // cos(160.3°)
        cos_table[115] = 31113;       // cos(161.7°)
        cos_table[116] = 31356;       // cos(163.1°)
        cos_table[117] = 31580;       // cos(164.5°)
        cos_table[118] = 31785;       // cos(165.9°)
        cos_table[119] = 31970;       // cos(167.3°)
        cos_table[120] = 32137;       // cos(168.8°)
        cos_table[121] = 32284;       // cos(170.2°)
        cos_table[122] = 32412;       // cos(171.6°)
        cos_table[123] = 32520;       // cos(173.0°)
        cos_table[124] = 32609;       // cos(174.4°)
        cos_table[125] = 32678;       // cos(175.8°)
        cos_table[126] = 32727;       // cos(177.2°)
        cos_table[127] = 32757;       // cos(178.6°)
    end
    logic [ANGLE_WIDTH-1:0] cos_angle;
    assign cos_angle = $unsigned(7'sd90 - angle);
    // Map input angle to LUT value

    assign sin_value = cos_table[cos_angle];
    assign sign_bit = cos_angle > 64;

endmodule

`default_nettype wire